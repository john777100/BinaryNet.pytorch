`define TEST_DATA_CNT 1
`define BIT_CNT 	8
`define CHANNEL_CNT	256
`define INPUT_DIM	10
`define OUTPUT_DIM	10
//`define KERNEL_SIZE 16
//`define RELU_THRESHOLD `KERNEL_SIZE/2

`define ACC_WIDTH 		32


`define FP_WIDTH 		8
`define FP_PARALLEL 	16
`define FP_MODEL_WIDTH 	784
`define FP_CLOCK 		40850


`define PRO_WIDTH 		2
`define PRO_CH_CNT		4
`define PRO_PARALLEL 	16
`define PRO_MODEL_WIDTH 784
`define PRO_CLOCK 		6.5

`define BIN_PARALLEL 	8
`define BIN_MODEL_WIDTH 784
`define BIN_CLOCK 		21611

